`define DATA_WIDTH 8
`define FIFO_WIDTH 4
`define FIFO_SIZE (1<<`FIFO_WIDTH)